`include "./defines.v"
`include "./memory_controller.v"
`include "./pc.v"

module if_stage (
    input clk,
    input rstn,
    input pause,

    output waiting
);

endmodule
